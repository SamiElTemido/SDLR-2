library IEEE;
use ieee.std_logic_1164.all;

entity SN74LS47	is
	port(
	CLK: in std_logic;
	RST: in std_logic;
	NIB: in std_logic_vector(3 downto 0);
	SEG: in std_logic_vecto(6 downto 0)
	);								   
end SN74LS47;

architecture Behavioral of SN74LS47 is
signal
begin 
end Behavioral;

